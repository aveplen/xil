`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:19:56 11/27/2022 
// Design Name: 
// Module Name:    fp_adder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fp_adder(
    input sign1,
    input sign2,
    input [3:0] exp1,
    input [3:0] exp2,
    input [7:0] frac1,
    input [7:0] frac2,
    input sign_out,
    input [3:0] exp_out,
    input [7:0] frac_out
    );


endmodule
